/*
  This module is used to send/receive string of ascii characters to/from the UART module
  - TX: The ascii string is formatted as follows: S:[temperature_high][temperature_low][humidity_high][humidity_low]\n
  - Rx: LEDs controlling format: L:[ascii_led_1][ascii_led_2]\n. e.g.: L:01\n (LED 1 ON, LED 2 OFF)
*/
module uart_string(
  input wire clk_100Mhz,
  input wire rst_n,

  input wire [7: 0] temperature,//data_heart_rate,
  input wire [7: 0] humidity,//data_spo2,

  input wire rx,
  output wire tx,

  output wire led_1,
  output wire led_2
);

  localparam [1:0] parity_type = 2'b01; // ODD parity
  localparam [1:0] baud_rate = 2'b10;   // 9600 baud
  // SEND_INTERVAL = Clock frequency (100 MHz) * Time (1 second) = 100,000,000 cycles
  localparam SEND_INTERVAL = 100_000_000; // 1 second

  wire tx_done, rx_done;

  reg [2:0] tx_index;  // Index for 8 characters
  reg [7:0] tx_data;
  reg send_start;
  reg [31:0] timer_count; // Timer counter for 1-second delay
  wire tx_busy;

  // ASCII message to send
  reg [6:0] tx_msg [0:7];

  integer temp;

  initial begin
    tx_msg[0] = 8'h53; // ASCII 'S'
    tx_msg[1] = 8'h3A; // ASCII ':'
    tx_msg[2] = 8'h30; // ASCII '0'
    tx_msg[3] = 8'h30; // ASCII '0'
    tx_msg[4] = 8'h30; // ASCII '0'
    tx_msg[5] = 8'h30; // ASCII '0'
    tx_msg[6] = 8'h0A; // ASCII '\n'
  end

  // Sending logic - TX Handler
  reg STATE_STR;
  always @(posedge clk_100Mhz or negedge rst_n) begin
    /*
      Handle the state machine for sending the string of ASCII characters every 1 second via UART
      You should control the SFM with 2 different clock domains: 100MHz and baud rate 9600
    */
    if (!rst_n) begin
      // Reset all states and signals
      tx_msg[0] <= 8'h53; // ASCII 'S'
      tx_msg[1] <= 8'h3A; // ASCII ':'
      tx_msg[2] <= 8'h30; // ASCII '0'
      tx_msg[3] <= 8'h30; // ASCII '0'
      tx_msg[4] <= 8'h30; // ASCII '0'
      tx_msg[5] <= 8'h30; // ASCII '0'
      tx_msg[6] <= 8'h0A; // ASCII '\n

      tx_index <= 0;
      send_start <= 0;
      timer_count <= 0;
      STATE_STR <= 0;
    end else begin
      case (STATE_STR)
        0: begin
          // Wait for 1-second interval
          if (timer_count == SEND_INTERVAL) begin
            timer_count <= 0;
            STATE_STR <= 1; // Transition to sending state
          end else begin
            timer_count <= timer_count + 1;
          end
        end
        1: begin
          // Update sensor data at the start of transmission
          if (tx_index == 0 && !tx_busy) begin
            tx_msg[2] <= temperature / 10 + 8'h30;
            tx_msg[3] <= temperature % 10 + 8'h30;
            tx_msg[4] <= humidity / 10 + 8'h30;
            tx_msg[5] <= humidity % 10 + 8'h30;
          end

          // Send one character at a time
          if (!tx_busy && !send_start) begin
            tx_data <= tx_msg[tx_index]; // Load the current character
            send_start <= 1;            // Start UART transmission
          end else if (!tx_busy && send_start) begin
            send_start <= 0;            // Clear send_start after transmission
            if (tx_index < 6) begin
              tx_index <= tx_index + 1; // Move to the next character
            end else begin
              tx_index <= 0;            // Reset index after all characters are sent
              STATE_STR <= 0;           // Transition back to idle state
            end
          end
        end
      endcase
    end
  end

  /*
  Rx Handler
  */
  reg [7:0] rx_msg [0:4]; // Buffer for received 5 characters
  reg [3:0] rx_index;  // Index for 4 characters
  wire [7:0] rx_data;
  reg led_1_reg, led_2_reg;
  assign led_1 = led_1_reg;
  assign led_2 = led_2_reg;
  wire rx_busy;
  always @(posedge clk_100Mhz or negedge rst_n) begin
    if (!rst_n) begin
      rx_index <= 0;
      
      rx_msg[0] <= 8'h4C; // ASCII 'L'
      rx_msg[1] <= 8'h3A; // ASCII ':'
      rx_msg[2] <= 8'h30; // ASCII '0'
      rx_msg[3] <= 8'h30; // ASCII '0'
      rx_msg[4] <= 8'h0A; // ASCII '\n'

      led_2_reg <= 1'b1;
      led_1_reg <= 1'b1;
    end else begin
      // if not busy and done receiving a character
      if (!rx_busy && rx_done) begin
        // ok, you have just received a character
        // let store it in the buffer
        rx_msg[rx_index] <= rx_data;

        // check if exceeds the buffer size:
        rx_index <= (rx_index < 4) ? rx_index + 1 : 0; // Increment or reset buffer index

        // check if it is a newline character (final character)
        if (rx_data == 8'h0A) begin
          rx_index <= 0;

          // done a string. e.g.: L:01\n
          // let control the LEDs
          if (rx_msg[0] == 8'h4C) begin // Check for 'L' (led)
            led_1_reg <= rx_msg[2] == 8'h31 ? 1'b1 : 1'b0;
            led_2_reg <= rx_msg[3] == 8'h31 ? 1'b1 : 1'b0;
          end
        end
      end else if (rx_done) begin
        led_2_reg <= 1'b0;
        led_1_reg <= 1'b0;
      end
    end
  end

  uart_tx uart_tx_inst(
    .clk(clk_100Mhz),
    .rst_n(rst_n),
    .tx_start(send_start),
    .tx_data(tx_data),
    .tx(tx),
    .tx_busy(tx_busy)
  );

  uart_rx uart_rx_inst (
    .clk(clk_100Mhz),
    .rst_n(rst_n),
    .rx(rx),
    .data_out(rx_data),
    .rx_busy(rx_busy),
    .done(rx_done)
  );
  /*
  TxUnit Transmitter(
    //  Inputs
    .reset_n(rst_n),
    .send(send_start),
    .clock(clk_100Mhz),
    .parity_type(parity_type),
    .baud_rate(baud_rate),
    .data_in(tx_data),

    //  Outputs
    .data_tx(tx),
    .active_flag(tx_busy),
    .done_flag(tx_done)
  );

  RxUnit Reciever(
    //  Inputs
    .reset_n(rst_n),
    .clock(clk_100Mhz),
    .parity_type(parity_type),
    .baud_rate(baud_rate),
    .data_tx(rx),

    //  Outputs
    .data_out(rx_data),
    .error_flag(),
    .active_flag(rx_busy),
    .done_flag(rx_done)
  );
  */

endmodule